`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Original file prepared by Mahdad Davari
// Modified and revised by Yuan Yao
//////////////////////////////////////////////////////////////////////////////////


module accelerator_tb # 
    (
        parameter integer INPUT_SIZE = 10,
        parameter integer RESULT_SIZE = 1,
        parameter integer WEIGHT_SIZE = INPUT_SIZE*RESULT_SIZE,
        parameter integer INPUT_ADDR_SIZE = 10, //[9:0]
        parameter integer RESULT_ADDR_SIZE = 2, //[5:0]
        parameter integer WEIGHT_ADDR_SIZE = 10, //[14:0]
        parameter integer FIXED_POINT_AMOUNT = 12, 
        parameter integer DATA_WIDTH = 32    
    )
    (

    );
    
    reg  s00_axi_aclk;
    reg  s00_axi_aresetn;

    // Ports of Axi Slave Bus Interface S00_AXIS
    wire  s00_axis_tready, valid_MAC_result;
    reg [DATA_WIDTH-1 : 0] s00_axis_tdata;
    reg [(DATA_WIDTH/8)-1 : 0] s00_axis_tstrb;
    reg  s00_axis_tlast;
    reg  s00_axis_tvalid;

    // Ports of Axi Master Bus Interface M00_AXIS
    wire  m00_axis_tvalid;
    wire [DATA_WIDTH-1 : 0] m00_axis_tdata, MAC_results;
    wire [(DATA_WIDTH/8)-1 : 0] m00_axis_tstrb;
    wire  m00_axis_tlast;
    reg  m00_axis_tready;
    
    reg sel;
    reg start;
    
    integer row;
    integer column;
    integer count;
    
    integer matRSW [0:RESULT_SIZE-1] = '{268};//, 119539, -38978, 12731, 37346}; //, 74829, 41561, -36134, -58525, -164845, 31255, -118765, -84873, -149139, -31484, 47832, -197099, 61694, 59350, -18467, 54140, -67870, 26591, -31328, 126714, -21026, 109507, -205420, -30868, 81067};
    integer matRHW [0:RESULT_SIZE-1];
    
  
	 


    
    integer image[0:INPUT_SIZE-1] = '{1, 1, 0, 0, 0, 0, 0, 0, 0, 0}; //, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1344, 2960, 2544, 2416, 960, 576, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3552, 4064, 4064, 4064, 4064, 3856, 3168, 3168, 3168, 3168, 3168, 3168, 3168, 3168, 2720, 832, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1072, 1824, 1152, 1824, 2608, 3632, 4064, 3600, 4064, 4064, 4064, 4000, 3664, 4064, 4064, 2240, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 272, 1056, 224, 1072, 1072, 1072, 944, 336, 3776, 4064, 1696, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1328, 4048, 3344, 288, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 352, 3728, 4080, 1328, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2064, 4064, 3808, 704, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 944, 3984, 4064, 992, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2128, 4064, 2992, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 144, 3280, 3968, 928, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2016, 4064, 2912, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1200, 4016, 3840, 912, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 304, 3536, 4064, 2656, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 3248, 4064, 3504, 560, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 608, 4064, 4064, 1232, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 496, 3584, 4064, 1840, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2128, 4064, 4064, 832, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 976, 3872, 4064, 4064, 832, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1936, 4064, 4064, 3504, 640, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1936, 4064, 3312, 288, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0}; 
    integer layer_0[0:WEIGHT_SIZE-1] = '{999999, 99999, -631, 6241, 2930, 1705, -7018, 207, -1440, 2801};// 4469, 1782, -1949, -568, 1367, -7916, -2099, 9340, 2955, -2352, -4583, 199, -3223, 3954, 6863, 157, -3506, -4008, -2747, -5039, 4486, -728, -3061, 9474, 2711, -781, 1190, -3427, -3313, -2769, -5597, -8668, 1857, -8920, -2868, -148, 2234, 798, -64, 1648, -626, -3606, 8547, 4212, -909, -2015, 539, 584, -1497, -3608, 3260, -1118, 1306, -5051, 6285, 2043, 2124, 6561, -6169, -2082, 5013, -4076, -570, -6644, -4191, -3264, 1701, -8820, 8626, -1448, 4714, 2082, -569, 3535, 4961, -3934, 1775, -6911, -2158, -2931, -353, 5851, -621, -2074, 2305, -2762, -613, 1279, 977, -12035, -3047, -4923, 1541, -1886, 3161, -2749, 5048, 5562, 5848, -3869, 1285, 909, -4251, 364, -3459, 2484, -3942, 3025, -1320, 3636, 1221, 7362, 5564, 4993, 1671, 11770, -2356, -6639, -828, -5173, 3039, -733, -238, -1628, 8591, -2101, -2692, -4723, 3402, -3841, -1682, 3864, 523, -2337, 2665, 2589, -62, -5378, -4509, 3637, 4508, 4108, 3789, -3442, -3338, -3942, 2065, 8287, 4349, 12487, 10055, 4585, 3339, 9006, 2029, 5517, 7056, 7344, 7194, -10241, -4092, 7779, -4840, -3673, 6467, 9491, -1778, -6426, 3531, 391, -6831, -69, 3825, -4401, -989, -446, -508, 1181, -1306, -2722, 4730, -3625, 311, 2662, 618, 6067, -2167, 1775, -643, -4871, 5092, 2358, -2959, 3575, 1772, -257, -9319, 2069, 2893, -5235, -4993, 1410, 4736, -5651, -8900, 1966, -4954, -516, 8871, 1557, 10314, -1356, -294, -1704, 1962, 1124, 1721, 3699, -5509, -8286, -4435, -7278, 830, 7209, -4211, -8481, 1277, -1155, -7056, 2522, -4305, 3518, -4550, 8330, -2366, 2777, -2865, 5825, 4349, 1024, 6292, 1115, -5110, 7287, 998, 3781, -3031, -3472, -8434, -3435, -7660, -3164, 2834, -780, -2090, -1228, 797, -3887, 185, -3971, -2135, -2618, -7515, -3377, -295, -1568, 10485, -2042, 4433, -9451, 3564, 4953, 2223, 842, 642, -4017, -3456, -2973, 2370, 871, -6863, -397, 491, -13164, -8986, -6708, -4440, -6588, -2558, -1397, -923, -5575, -4310, -2206, 2506, 4927, -916, 5155, -447, 1400, -964, 1365, -3584, 10815, -2214, 306, 2618, 4200, 2172, 546, -1011, -3270, -12047, -7912, 265, 4408, 757, -5490, -1301, -2254, 5392, 8977, 2329, -263, -1275, 242, 3245, -917, 4890, 1068, -1580, -1279, 7981, -4960, -1687, -3945, 3292, 2140, 7941, -4580, 4216, 2302, -3214, -944, 475, 4019, 977, -655, -2478, 4876, -3101, -3467, -5021, -1641, 1444, -2744, -6311, -1229, -1658, 594, 4037, -580, 161, 7884, 4708, 5475, 14245, 18296, 3281, 3043, -2904, -3428, 4374, 3193, 3124, 4428, 6196, 4094, -4547, -486, 4872, 4442, -2312, 6599, 843, 6036, 931, 5417, -3071, 10201, 6593, 3025, 537, 7310, 19539, 9788, 990, 428, 3476, 3760, -6816, -726, -4125, 9905, -2572, 3377, -5495, 2760, -613, -429, -352, -3041, -782, -1350, -581, 6312, 2159, 3264, 4487, -5162, 551, 13338, 12167, 2006, -9677, 13231, 135, -198, -7276, -10774, -2546, -7653, -4763, 9057, -3133, 2055, -1297, -3774, -7281, 10980, 3123, 1920, -5667, 3245, 5291, -7014, 1752, 3361, 8237, 19829, 4571, 210, 2752, 2533, -2142, 3036, 2279, -817, -9290, -1975, -5906, -1462, 2096, 1342, -352, -237, 5855, 202, -2019, 1877, -4593, 7607, 9203, 1, 1826, 5665, 9883, 13423, 2813, -1183, -8729, -2269, 531, -4886, -3083, -4765, -4602, 1769, -3776, 3920, -1526, -1324, -1210, 39, 1384, 2415, 1845, 4969, -978, -5661, 8928, -3340, 6071, 12403, 4760, 10001, -542, -9803, -1419, 2432, 5239, -2958, -6537, 1950, 1584, 3901, -1042, 2005, 7866, -1420, -5519, 3312, 2338, 1303, -3478, 5735, -1414, 4752, 8851, 1108, 11302, 5608, -4334, 7674, 1462, 1066, -11, -2282, -3207, 6636, 3373, 3037, 7477, 4559, 1017, -1426, 7787, 6486, -1612, 3303, 10824, 3321, -3383, 1822, -4878, 4088, 7536, 3668, 7146, 2175, 10291, 1349, 3631, -1798, -4770, -6639, 2905, 2883, 7998, 2122, 10099, 13353, 6589, 1502, 1402, -3743, 730, -2639, 1998, 2781, 7971, 1071, 4650, 8399, 7245, 4807, -2393, 1510, -90, 1390, 1821, 257, 1379, -1035, 1969, 5976, 5553, 4870, 7174, 6831, 8142, 3466, -2632, 6040, -7988, 3290, 2772, 3069, -1191, 709, 4001, 7714, 835, 647, 2816, -8212, 8931, -853, -928, 1344, -1753, 4545, -447, -1995, 7303, 230, 10218, 3896, -1055, 1477, 7548, 98, -3255, -2023, 1828, 4389, 729, 5015, -9300, -3374, -5469, -13483, -643, 4017, 7198, 637, 8457, 464, -430, 1982, -1300, -1716, -3750, 9128, 110, -681, 2497, 2743, -1339, 1598, -1359, 218, 5695, 108, 1226, -3672, -6679, 157, -6371, -3495, -3528, -3958, 4145, 1536, -3526, -3892, 3173, 6458, 6525, 174, 4682, -2040, -4541, 4103, 1289, 521, 1908, -95, 1520, -5236, -1103, 7658, 1568, -3085, 559, 6608, 4142, -9729, -1951, -5576, -3926, -1208, -945, 1656, 718, -3001, -589, -1237, 3946, 4614, 1176, 983, -3266, 8166, -558, -6957, -5895, -6724, -6085, 2315, 1863, -2157, -438, 5584, 1240, 766, -3500, 1252, 5196, -6853, 1299, 4427, 1364, 539, 4460, -451, -1940, 1781, -1204, -3897, -3166, -689, -2021, -2902, 3669, -2803, -6068, 4829, -3160, 3303, 2230, 759, 65, -1865, 3389, 416, 1340, 488, -854, -3584, 363, -5876, -2125, 3222, -1718, -3476, 5565, 4193, -1150, -601, -7274, 1159, 4700, -4627};


    
    mat_mul # (
    .INPUT_SIZE(INPUT_SIZE),
    .RESULT_SIZE (RESULT_SIZE),
    .WEIGHT_SIZE (WEIGHT_SIZE),
    .INPUT_ADDR_SIZE(INPUT_ADDR_SIZE),
    .RESULT_ADDR_SIZE(RESULT_ADDR_SIZE),
    .WEIGHT_ADDR_SIZE(WEIGHT_ADDR_SIZE),
    .FIXED_POINT_AMOUNT(FIXED_POINT_AMOUNT),
    .DATA_WIDTH(DATA_WIDTH)    
    ) accelerator (
    .s00_axi_aclk(s00_axi_aclk),
    .s00_axi_aresetn(s00_axi_aresetn),
    .s00_axis_tready(s00_axis_tready),
    .s00_axis_tdata(s00_axis_tdata),
    .s00_axis_tlast(s00_axis_tlast),
    .s00_axis_tvalid(s00_axis_tvalid),
    .m00_axis_tvalid(m00_axis_tvalid),
    .m00_axis_tdata(m00_axis_tdata),
    .m00_axis_tstrb(m00_axis_tstrb),
    .m00_axis_tlast(m00_axis_tlast),
    .m00_axis_tready(m00_axis_tready),
    .sel(sel),
    .start(start),
    .MAC_result(MAC_results),
    .valid_MAC_result(valid_MAC_result)
    );
    wire temporary_permanent_value;
    reg [DATA_WIDTH-1 : 0] slv_reg1;
    reg permanent_valid;
    always @ (valid_MAC_result, MAC_results, temporary_permanent_value) begin
        if (valid_MAC_result) begin
            slv_reg1 = MAC_results;
            permanent_valid <= 1; end
    end
    
    
    always
        #10 s00_axi_aclk = ~s00_axi_aclk;
        
    initial begin
        s00_axi_aclk = 1;
        s00_axi_aresetn = 0;
        s00_axis_tdata = 0;
        s00_axis_tstrb = 4'hf;
        s00_axis_tlast = 0;
        s00_axis_tvalid = 0;
        m00_axis_tready = 0;
        sel = 0;
        start = 0;
        row = 0;
        column = 0;
        count = 0;
        
        // initialise the matrices; for debug use $urandom%10 to have unsigned values less than 10;
        // $srandom(12345); // Uncomment for debug, which will always generates the same random numbers
        for (row = 0; row < RESULT_SIZE; row = row + 1) begin
                matRHW [row] = 0;
        end
        
        
        #20
        s00_axi_aresetn = 1;
        count = 0;
        
        // send the two matrices using the AXI Stream protocol
        $display ("LOADING WEIGHTS");
        #20
        s00_axis_tvalid = 1;
        for (row = 0; row < WEIGHT_SIZE; row = row + 1) begin
                // Should use non-blocking assignment here
                s00_axis_tdata <= layer_0[row];
                
                // set the last signal when sending the last data item
                if (row == WEIGHT_SIZE-1)
                    s00_axis_tlast = 1;
                #20;
                
                // wait until the slave is ready to read the data
                while (!s00_axis_tready) begin
                    #20;
                end
        end
        
        s00_axis_tlast = 0;
        s00_axis_tvalid = 0;
        
        
        //SEND INPUT
        $display ("LOADING IMAGE");
        sel = 1;

        #20
        s00_axi_aresetn = 1;
        count = 0;
        
        // send the two matrices using the AXI Stream protocol
        #20
        s00_axis_tvalid = 1;
        for (row = 0; row < INPUT_SIZE; row = row + 1) begin
            // Should use non-blocking assignment here
            s00_axis_tdata <= image[row];
            
            // set the last signal when sending the last data item
            if (row == INPUT_SIZE-1)
                s00_axis_tlast = 1;
            #20;
            
            // wait until the slave is ready to read the data
            while (!s00_axis_tready) begin
                #20;
            end
        end
        
        s00_axis_tlast = 0;
        s00_axis_tvalid = 0;
        
        
        // START the accelerator
        $display ("STARTING ACCELERATOR");
        #20
        start = 1;
        #20
        start = 0;
        
        // wait for the reslt to arrive from the accelerator
        m00_axis_tready = 1;
        
        row = 0;
        $display("WAITING FOR ACCELERATOR TO FINISH");
        while (!m00_axis_tlast) begin // exit if last data already received
            #20;
            if (m00_axis_tvalid == 1) begin // valid data on the bus
                matRHW[row] = m00_axis_tdata;
                row = row + 1;
            end
        end
        $display("GETTING RESULT");
        
        m00_axis_tready = 0;
        count = 0;
        $display("COMPARING RESULT");
        // compare the hardware and software results
        for (row = 0; row < RESULT_SIZE; row = row + 1) begin
            $display("%d", matRHW[row]);
            $display("ROW %d", row);
            if (matRSW [row] != matRHW [row] || ^matRHW [row] === 1'bX) begin
                count = count + 1;
                $display ("HW/SW result mismatch! row=%d; res_sw=%d; res_hw=%d", row, matRSW[row], matRHW[row]);
            end
        end

       if (count == 0)
            $display ("HW/SW result match!");
       #40
       $stop;
       
    end
    
endmodule